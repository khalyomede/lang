module lang

pub fn Lang.from_iso_2(code string) ?Lang {
    return match code {
        'aa' { Lang.aa }
        'ab' { Lang.ab }
        'af' { Lang.af }
        'ak' { Lang.ak }
        'sq' { Lang.sq }
        'am' { Lang.am }
        'ar' { Lang.ar }
        'an' { Lang.an }
        'hy' { Lang.hy }
        'as' { Lang.as }
        'av' { Lang.av }
        'ae' { Lang.ae }
        'ay' { Lang.ay }
        'az' { Lang.az }
        'ba' { Lang.ba }
        'bm' { Lang.bm }
        'eu' { Lang.eu }
        'be' { Lang.be }
        'bn' { Lang.bn }
        'bi' { Lang.bi }
        'bo' { Lang.bo }
        'bs' { Lang.bs }
        'br' { Lang.br }
        'bg' { Lang.bg }
        'my' { Lang.my }
        'ca' { Lang.ca }
        'ch' { Lang.ch }
        'ce' { Lang.ce }
        'zh' { Lang.zh }
        'cu' { Lang.cu }
        'cv' { Lang.cv }
        'kw' { Lang.kw }
        'co' { Lang.co }
        'cr' { Lang.cr }
        'cs' { Lang.cs }
        'da' { Lang.da }
        'dv' { Lang.dv }
        'nl' { Lang.nl }
        'dz' { Lang.dz }
        'en' { Lang.en }
        'eo' { Lang.eo }
        'et' { Lang.et }
        'ee' { Lang.ee }
        'fo' { Lang.fo }
        'fa' { Lang.fa }
        'fj' { Lang.fj }
        'fi' { Lang.fi }
        'fr' { Lang.fr }
        'ff' { Lang.ff }
        'fy' { Lang.fy }
        'gd' { Lang.gd }
        'ga' { Lang.ga }
        'gl' { Lang.gl }
        'gv' { Lang.gv }
        'el' { Lang.el }
        'gn' { Lang.gn }
        'gu' { Lang.gu }
        'ht' { Lang.ht }
        'ha' { Lang.ha }
        'he' { Lang.he }
        'hz' { Lang.hz }
        'hi' { Lang.hi }
        'ho' { Lang.ho }
        'hr' { Lang.hr }
        'hu' { Lang.hu }
        'ig' { Lang.ig }
        'is' { Lang.is }
        'io' { Lang.io }
        'ii' { Lang.ii }
        'iu' { Lang.iu }
        'ie' { Lang.ie }
        'ia' { Lang.ia }
        'id' { Lang.id }
        'ik' { Lang.ik }
        'it' { Lang.it }
        'jv' { Lang.jv }
        'ja' { Lang.ja }
        'kl' { Lang.kl }
        'kn' { Lang.kn }
        'ks' { Lang.ks }
        'ka' { Lang.ka }
        'kr' { Lang.kr }
        'kk' { Lang.kk }
        'km' { Lang.km }
        'ki' { Lang.ki }
        'rw' { Lang.rw }
        'ky' { Lang.ky }
        'kv' { Lang.kv }
        'kg' { Lang.kg }
        'ko' { Lang.ko }
        'kj' { Lang.kj }
        'ku' { Lang.ku }
        'lo' { Lang.lo }
        'la' { Lang.la }
        'lv' { Lang.lv }
        'li' { Lang.li }
        'ln' { Lang.ln }
        'lt' { Lang.lt }
        'lb' { Lang.lb }
        'lu' { Lang.lu }
        'lg' { Lang.lg }
        'mk' { Lang.mk }
        'mh' { Lang.mh }
        'ml' { Lang.ml }
        'mi' { Lang.mi }
        'mr' { Lang.mr }
        'ms' { Lang.ms }
        'mg' { Lang.mg }
        'mt' { Lang.mt }
        'mn' { Lang.mn }
        'na' { Lang.na }
        'nv' { Lang.nv }
        'nr' { Lang.nr }
        'nd' { Lang.nd }
        'ng' { Lang.ng }
        'ne' { Lang.ne }
        'nn' { Lang.nn }
        'nb' { Lang.nb }
        'no' { Lang.no }
        'ny' { Lang.ny }
        'oc' { Lang.oc }
        'oj' { Lang.oj }
        'or' { Lang.or }
        'om' { Lang.om }
        'os' { Lang.os }
        'pa' { Lang.pa }
        'pi' { Lang.pi }
        'pl' { Lang.pl }
        'pt' { Lang.pt }
        'ps' { Lang.ps }
        'qu' { Lang.qu }
        'rm' { Lang.rm }
        'ro' { Lang.ro }
        'rn' { Lang.rn }
        'ru' { Lang.ru }
        'sg' { Lang.sg }
        'sa' { Lang.sa }
        'si' { Lang.si }
        'sk' { Lang.sk }
        'sl' { Lang.sl }
        'se' { Lang.se }
        'sm' { Lang.sm }
        'sn' { Lang.sn }
        'sd' { Lang.sd }
        'so' { Lang.so }
        'st' { Lang.st }
        'es' { Lang.es }
        'sc' { Lang.sc }
        'sr' { Lang.sr }
        'ss' { Lang.ss }
        'su' { Lang.su }
        'sw' { Lang.sw }
        'sv' { Lang.sv }
        'ty' { Lang.ty }
        'ta' { Lang.ta }
        'tt' { Lang.tt }
        'te' { Lang.te }
        'tg' { Lang.tg }
        'tl' { Lang.tl }
        'th' { Lang.th }
        'ti' { Lang.ti }
        'to' { Lang.to }
        'tn' { Lang.tn }
        'ts' { Lang.ts }
        'tk' { Lang.tk }
        'tr' { Lang.tr }
        'tw' { Lang.tw }
        'ug' { Lang.ug }
        'uk' { Lang.uk }
        'ur' { Lang.ur }
        'uz' { Lang.uz }
        've' { Lang.ve }
        'vi' { Lang.vi }
        'vo' { Lang.vo }
        'cy' { Lang.cy }
        'wa' { Lang.wa }
        'wo' { Lang.wo }
        'xh' { Lang.xh }
        'yi' { Lang.yi }
        'yo' { Lang.yo }
        'za' { Lang.za }
        'zu' { Lang.zu }
        else { none }
    }
}
